module api

import interfaces

pub fn Window.new() interfaces.Window {
	return Window{}
}