module unbreakable

pub struct Sprite {
	GameObject
}
