module unbreakable

// pub interface Renderable {
// }

struct DrawManager {
	geometry Geometry
}

fn (self DrawManager) render() {
}

fn init_draw_manager() DrawManager {
	return DrawManager{}
}
