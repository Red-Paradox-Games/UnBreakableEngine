module unbreakable

struct Geometry {
}
