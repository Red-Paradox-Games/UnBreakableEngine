module unbreakable