module unbreakable

fn main() {
	println('Hello World!')
}
