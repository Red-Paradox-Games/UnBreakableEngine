module graphics
